"","Phase","Item.Type","Block","Item.Number","Talker.A","Talker.A_Materials","Talker.A_Sound","Talker.B","Talker.B_Materials","Talker.B_Sound","Version","Talker.A_Gender","Talker.A_Ear","Talker.B_Gender","Talker.B_Ear","rep","filename"
"1","Exposure","Critical",1,1,"Ambition","Materials A","Sh","Parasite","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Ambition.M.L_NAS.Parasite.F.R.wav"
"2","Exposure","Critical",1,2,"Machinery","Materials A","Sh","Obscene","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Machinery.M.L_NAS.Obscene.F.R.wav"
"3","Exposure","Critical",1,3,"Brochure","Materials A","Sh","Medicine","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Brochure.M.L_NAS.Medicine.F.R.wav"
"4","Exposure","Critical",1,4,"Official","Materials A","Sh","Tennessee","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Official.M.L_NAS.Tennessee.F.R.wav"
"5","Exposure","Critical",1,5,"Crucial","Materials A","Sh","Penninsula","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Crucial.M.L_NAS.Penninsula.F.R.wav"
"6","Exposure","Critical",1,6,"Pediatrician","Materials A","Sh","Hallucinate","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Pediatrician.M.L_NAS.Hallucinate.F.R.wav"
"7","Exposure","Critical",1,7,"Flourishing","Materials A","Sh","Arkansas","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Flourishing.M.L_NAS.Arkansas.F.R.wav"
"8","Exposure","Critical",1,8,"Reassure","Materials A","Sh","Compensate","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Reassure.M.L_NAS.Compensate.F.R.wav"
"9","Exposure","Critical",1,9,"Graduation","Materials A","Sh","Dinosaur","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Graduation.M.L_NAS.Dinosaur.F.R.wav"
"10","Exposure","Critical",1,10,"Vacation","Materials A","Sh","Rehearsal","Materials B","S","Unshifted","Male","Left","Female","Right",1,"Critical_07.A_Sh.Vacation.M.L_NAS.Rehearsal.F.R.wav"
"11","Exposure","Critical",1,11,"Pregnancy","Materials B","S","Initial","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Pregnancy.M.L_A_Ash.Initial.F.R.wav"
"12","Exposure","Critical",1,12,"Democracy","Materials B","S","Beneficial","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Democracy.M.L_A_Ash.Beneficial.F.R.wav"
"13","Exposure","Critical",1,13,"Embassy","Materials B","S","Negotiate","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Embassy.M.L_A_Ash.Negotiate.F.R.wav"
"14","Exposure","Critical",1,14,"Legacy","Materials B","S","Commercial","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Legacy.M.L_A_Ash.Commercial.F.R.wav"
"15","Exposure","Critical",1,15,"Reconcile","Materials B","S","Parachute","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Reconcile.M.L_A_Ash.Parachute.F.R.wav"
"16","Exposure","Critical",1,16,"Personal","Materials B","S","Efficient","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Personal.M.L_A_Ash.Efficient.F.R.wav"
"17","Exposure","Critical",1,17,"Eraser","Materials B","S","Publisher","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Eraser.M.L_A_Ash.Publisher.F.R.wav"
"18","Exposure","Critical",1,18,"Episode","Materials B","S","Glacier","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Episode.M.L_A_Ash.Glacier.F.R.wav"
"19","Exposure","Critical",1,19,"Literacy","Materials B","S","Refreshing","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Literacy.M.L_A_Ash.Refreshing.F.R.wav"
"20","Exposure","Critical",1,20,"Coliseum","Materials B","S","Impatient","Materials A","Sh","Shifted","Male","Left","Female","Right",1,"Critical_07.B_As.Coliseum.M.L_A_Ash.Impatient.F.R.wav"
"21","Exposure","Filler",1,1,"America","Set A","Word","Wominid","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.America.F.R_N.Wominid.M.L.wav"
"22","Exposure","Filler",1,1,"Bakery","Set B","Word","Wojalto","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Bakery.M.L_N.Wojalto.F.R.wav"
"23","Exposure","Filler",1,1,"Ballerina","Set C","Word","Youmgel","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Ballerina.M.R_N.Youmgel.F.L.wav"
"24","Exposure","Filler",1,2,"Blueberry","Set A","Word","Ungelnin","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Blueberry.F.R_N.Ungelnin.M.L.wav"
"25","Exposure","Filler",1,2,"Bullying","Set B","Word","Tounamplem","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Bullying.M.L_N.Tounamplem.F.R.wav"
"26","Exposure","Filler",1,2,"Burglary","Set C","Word","Tymolape","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Burglary.M.R_N.Tymolape.F.L.wav"
"27","Exposure","Filler",1,3,"Camera","Set A","Word","Tilegkalo","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Camera.F.R_N.Tilegkalo.M.L.wav"
"28","Exposure","Filler",1,3,"Continually","Set B","Word","Ryligal","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Continually.M.L_N.Ryligal.F.R.wav"
"29","Exposure","Filler",1,3,"Domineering","Set C","Word","Tamical","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Domineering.M.R_N.Tamical.F.L.wav"
"30","Exposure","Filler",1,4,"Directory","Set A","Word","Rimkeluwar","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Directory.F.R_N.Rimkeluwar.M.L.wav"
"31","Exposure","Filler",1,4,"Document","Set B","Word","Rawamtee","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Document.M.L_N.Rawamtee.F.R.wav"
"32","Exposure","Filler",1,4,"Embody","Set C","Word","Rengime","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Embody.M.R_N.Rengime.F.L.wav"
"33","Exposure","Filler",1,5,"Dynamite","Set A","Word","Rakil","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Dynamite.F.R_N.Rakil.M.L.wav"
"34","Exposure","Filler",1,5,"Eighty","Set B","Word","Ploupelai","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Eighty.M.L_N.Ploupelai.F.R.wav"
"35","Exposure","Filler",1,5,"Gullible","Set C","Word","Pourilar","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Gullible.M.R_N.Pourilar.F.L.wav"
"36","Exposure","Filler",1,6,"Gardenia","Set A","Word","Perkum","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Gardenia.F.R_N.Perkum.M.L.wav"
"37","Exposure","Filler",1,6,"Grammatical","Set B","Word","Omperoge","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Grammatical.M.L_N.Omperoge.F.R.wav"
"38","Exposure","Filler",1,6,"Honeymoon","Set C","Word","Almikquary","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Honeymoon.M.R_N.Almikquary.F.L.wav"
"39","Exposure","Filler",1,7,"Hamburger","Set A","Word","Nomerae","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Hamburger.F.R_N.Nomerae.M.L.wav"
"40","Exposure","Filler",1,7,"Identical","Set B","Word","Nempring","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Identical.M.L_N.Nempring.F.R.wav"
"41","Exposure","Filler",1,7,"Illuminate","Set C","Word","Niritaly","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Illuminate.M.R_N.Niritaly.F.L.wav"
"42","Exposure","Filler",1,8,"Hurdle","Set A","Word","Namuary","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Hurdle.F.R_N.Namuary.M.L.wav"
"43","Exposure","Filler",1,8,"Interior","Set B","Word","Mibgem","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Interior.M.L_N.Mibgem.F.R.wav"
"44","Exposure","Filler",1,8,"Ironic","Set C","Word","Makid","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Ironic.M.R_N.Makid.F.L.wav"
"45","Exposure","Filler",1,9,"Inhabit","Set A","Word","Logelai","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Inhabit.F.R_N.Logelai.M.L.wav"
"46","Exposure","Filler",1,9,"Knowingly","Set B","Word","Meidnow","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Knowingly.M.L_N.Meidnow.F.R.wav"
"47","Exposure","Filler",1,9,"Laminate","Set C","Word","Kaldemia","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Laminate.M.R_N.Kaldemia.F.L.wav"
"48","Exposure","Filler",1,10,"Keyboard","Set A","Word","Lenediaw","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Keyboard.F.R_N.Lenediaw.M.L.wav"
"49","Exposure","Filler",1,10,"Lethal","Set B","Word","Kermimer","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Lethal.M.L_N.Kermimer.F.R.wav"
"50","Exposure","Filler",1,10,"Liability","Set C","Word","Imdalier","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Liability.M.R_N.Imdalier.F.L.wav"
"51","Exposure","Filler",1,11,"Lengthen","Set A","Word","Kelabidel","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Lengthen.F.R_N.Kelabidel.M.L.wav"
"52","Exposure","Filler",1,11,"Lobbying","Set B","Word","Itempider","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Lobbying.M.L_N.Itempider.F.R.wav"
"53","Exposure","Filler",1,11,"Marina","Set C","Word","Kloumidiger","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Marina.M.R_N.Kloumidiger.F.L.wav"
"54","Exposure","Filler",1,12,"Lingering","Set A","Word","Inpaki","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Lingering.F.R_N.Inpaki.M.L.wav"
"55","Exposure","Filler",1,12,"Membrane","Set B","Word","Aknid","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Membrane.M.L_N.Aknid.F.R.wav"
"56","Exposure","Filler",1,12,"Metrical","Set C","Word","Halomimoc","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Metrical.M.R_N.Halomimoc.F.L.wav"
"57","Exposure","Filler",1,13,"Melancholy","Set A","Word","Hintarber","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Melancholy.F.R_N.Hintarber.M.L.wav"
"58","Exposure","Filler",1,13,"Negate","Set B","Word","Ibirak","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Negate.M.L_N.Ibirak.F.R.wav"
"59","Exposure","Filler",1,13,"Nightmare","Set C","Word","Gerbualo","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Nightmare.M.R_N.Gerbualo.F.L.wav"
"60","Exposure","Filler",1,14,"Napkin","Set A","Word","Gardimuallay","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Napkin.F.R_N.Gardimuallay.M.L.wav"
"61","Exposure","Filler",1,14,"Outnumber","Set B","Word","Halken","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Outnumber.M.L_N.Halken.F.R.wav"
"62","Exposure","Filler",1,14,"Panicking","Set C","Word","Galliwinou","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Panicking.M.R_N.Galliwinou.F.L.wav"
"63","Exposure","Filler",1,15,"Ornament","Set A","Word","Gairelom","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Ornament.F.R_N.Gairelom.M.L.wav"
"64","Exposure","Filler",1,15,"Parakeet","Set B","Word","Ganla","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Parakeet.M.L_N.Ganla.F.R.wav"
"65","Exposure","Filler",1,15,"Pilgrim","Set C","Word","Emhoutic","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Pilgrim.M.R_N.Emhoutic.F.L.wav"
"66","Exposure","Filler",1,16,"Pineapple","Set A","Word","Bikanian","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Pineapple.F.R_N.Bikanian.M.L.wav"
"67","Exposure","Filler",1,16,"Platonic","Set B","Word","Dadigal","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Platonic.M.L_N.Dadigal.F.R.wav"
"68","Exposure","Filler",1,16,"Predict","Set C","Word","Dilkuaund","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Predict.M.R_N.Dilkuaund.F.L.wav"
"69","Exposure","Filler",1,17,"Purgatory","Set A","Word","Baliber","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Purgatory.F.R_N.Baliber.M.L.wav"
"70","Exposure","Filler",1,17,"Tactical","Set B","Word","Bamtell","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Tactical.M.L_N.Bamtell.F.R.wav"
"71","Exposure","Filler",1,17,"Terminal","Set C","Word","Bowidai","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Terminal.M.R_N.Bowidai.F.L.wav"
"72","Exposure","Filler",1,18,"Therapeutic","Set A","Word","Amalar","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Therapeutic.F.R_N.Amalar.M.L.wav"
"73","Exposure","Filler",1,18,"Titanium","Set B","Word","Anemer","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Titanium.M.L_N.Anemer.F.R.wav"
"74","Exposure","Filler",1,18,"Turbulent","Set C","Word","Anolipa","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Turbulent.M.R_N.Anolipa.F.L.wav"
"75","Exposure","Filler",1,19,"Tutorial","Set A","Word","Ailounam","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Tutorial.F.R_N.Ailounam.M.L.wav"
"76","Exposure","Filler",1,19,"Umbrella","Set B","Word","Lilgrai","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Umbrella.M.L_N.Lilgrai.F.R.wav"
"77","Exposure","Filler",1,19,"Undermine","Set C","Word","Alnadiro","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Undermine.M.R_N.Alnadiro.F.L.wav"
"78","Exposure","Filler",1,20,"Wealthy","Set A","Word","Acomining","Set A","Nonword","3","Female","Right","Male","Left",1,"Filler_A.03_W.Wealthy.F.R_N.Acomining.M.L.wav"
"79","Exposure","Filler",1,20,"Worldly","Set B","Word","Admunker","Set B","Nonword","4","Male","Left","Female","Right",1,"Filler_B.04_W.Worldly.M.L_N.Admunker.F.R.wav"
"80","Exposure","Filler",1,20,"Wrinkle","Set C","Word","Aigi","Set C","Nonword","1","Male","Right","Female","Left",1,"Filler_C.01_W.Wrinkle.M.R_N.Aigi.F.L.wav"
"81","Test","Test",3,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.03_F.1.ashi.25.wav"
"82","Test","Test",4,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.04_F.1.ashi.25.wav"
"83","Test","Test",7,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.07_F.1.ashi.25.wav"
"84","Test","Test",8,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.08_F.1.ashi.25.wav"
"85","Test","Test",11,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.11_F.1.ashi.25.wav"
"86","Test","Test",12,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.12_F.1.ashi.25.wav"
"87","Test","Test",1,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.01_M.1.ashi.25.wav"
"88","Test","Test",2,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.02_M.1.ashi.25.wav"
"89","Test","Test",5,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.05_M.1.ashi.25.wav"
"90","Test","Test",6,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.06_M.1.ashi.25.wav"
"91","Test","Test",9,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.09_M.1.ashi.25.wav"
"92","Test","Test",10,1,"ashi.25",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.10_M.1.ashi.25.wav"
"93","Test","Test",3,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.03_F.2.ashi.30.wav"
"94","Test","Test",4,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.04_F.2.ashi.30.wav"
"95","Test","Test",7,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.07_F.2.ashi.30.wav"
"96","Test","Test",8,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.08_F.2.ashi.30.wav"
"97","Test","Test",11,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.11_F.2.ashi.30.wav"
"98","Test","Test",12,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.12_F.2.ashi.30.wav"
"99","Test","Test",1,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.01_M.2.ashi.30.wav"
"100","Test","Test",2,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.02_M.2.ashi.30.wav"
"101","Test","Test",5,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.05_M.2.ashi.30.wav"
"102","Test","Test",6,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.06_M.2.ashi.30.wav"
"103","Test","Test",9,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.09_M.2.ashi.30.wav"
"104","Test","Test",10,2,"ashi.30",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.10_M.2.ashi.30.wav"
"105","Test","Test",3,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.03_F.3.ashi.40.wav"
"106","Test","Test",4,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.04_F.3.ashi.40.wav"
"107","Test","Test",7,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.07_F.3.ashi.40.wav"
"108","Test","Test",8,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.08_F.3.ashi.40.wav"
"109","Test","Test",11,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.11_F.3.ashi.40.wav"
"110","Test","Test",12,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.12_F.3.ashi.40.wav"
"111","Test","Test",1,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.01_M.3.ashi.40.wav"
"112","Test","Test",2,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.02_M.3.ashi.40.wav"
"113","Test","Test",5,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.05_M.3.ashi.40.wav"
"114","Test","Test",6,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.06_M.3.ashi.40.wav"
"115","Test","Test",9,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.09_M.3.ashi.40.wav"
"116","Test","Test",10,3,"ashi.40",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.10_M.3.ashi.40.wav"
"117","Test","Test",3,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.03_F.4.ashi.45.wav"
"118","Test","Test",4,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.04_F.4.ashi.45.wav"
"119","Test","Test",7,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.07_F.4.ashi.45.wav"
"120","Test","Test",8,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.08_F.4.ashi.45.wav"
"121","Test","Test",11,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.11_F.4.ashi.45.wav"
"122","Test","Test",12,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.12_F.4.ashi.45.wav"
"123","Test","Test",1,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.01_M.4.ashi.45.wav"
"124","Test","Test",2,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.02_M.4.ashi.45.wav"
"125","Test","Test",5,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.05_M.4.ashi.45.wav"
"126","Test","Test",6,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.06_M.4.ashi.45.wav"
"127","Test","Test",9,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.09_M.4.ashi.45.wav"
"128","Test","Test",10,4,"ashi.45",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.10_M.4.ashi.45.wav"
"129","Test","Test",3,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.03_F.5.ashi.50.wav"
"130","Test","Test",4,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.04_F.5.ashi.50.wav"
"131","Test","Test",7,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.07_F.5.ashi.50.wav"
"132","Test","Test",8,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.08_F.5.ashi.50.wav"
"133","Test","Test",11,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.11_F.5.ashi.50.wav"
"134","Test","Test",12,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.12_F.5.ashi.50.wav"
"135","Test","Test",1,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.01_M.5.ashi.50.wav"
"136","Test","Test",2,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.02_M.5.ashi.50.wav"
"137","Test","Test",5,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.05_M.5.ashi.50.wav"
"138","Test","Test",6,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.06_M.5.ashi.50.wav"
"139","Test","Test",9,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.09_M.5.ashi.50.wav"
"140","Test","Test",10,5,"ashi.50",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.10_M.5.ashi.50.wav"
"141","Test","Test",3,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.03_F.6.ashi.70.wav"
"142","Test","Test",4,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.04_F.6.ashi.70.wav"
"143","Test","Test",7,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.07_F.6.ashi.70.wav"
"144","Test","Test",8,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.08_F.6.ashi.70.wav"
"145","Test","Test",11,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.11_F.6.ashi.70.wav"
"146","Test","Test",12,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Female",NA,NA,NA,1,"Test_B.12_F.6.ashi.70.wav"
"147","Test","Test",1,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.01_M.6.ashi.70.wav"
"148","Test","Test",2,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.02_M.6.ashi.70.wav"
"149","Test","Test",5,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.05_M.6.ashi.70.wav"
"150","Test","Test",6,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.06_M.6.ashi.70.wav"
"151","Test","Test",9,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.09_M.6.ashi.70.wav"
"152","Test","Test",10,6,"ashi.70",NA,NA,NA,NA,NA,NA,"Male",NA,NA,NA,1,"Test_B.10_M.6.ashi.70.wav"
